package decode_test_pkg;
  
  import uvm_pkg::*;
  import uvmf_base_pkg::*;
  import lc3_env_pkg::*;
  
  `include "uvm_macros.svh"

  `include "lc3_test_pkg/test_top.sv"

endpackage